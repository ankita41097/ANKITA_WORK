jxjshxushsu
