module test;

input a;        
input b;

my name is ankita banerjee
$display(single line comment should be removed);
endmoduleinput a;
$display(single line comment should be removed);
