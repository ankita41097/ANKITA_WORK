module test;
/* This is multi line comment
it should be removed*/
input a;        //inline comment should be removed
input b;
//$display("a,b\n");//$display(single line comment should be removed);
/*$display(single line comment should be removed)*/my name is ankita banerjee//my name is;$displayjghjfhjfh
$display(single line comment should be removed);
endmodule/*$display(single line comment should be removed);*/input a;//$display(single line comment should be removed);
$display(single line comment should be removed);
