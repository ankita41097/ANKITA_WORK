module test;
input a;
input b;//inline comments//display("my name is ankita");/*this is multi line comment should be removed*/
$display("this is display statement");
$display();input b;//inline comments//display("my name is ankita");/*this is multi line comment should be removed*/
input b;//inline comments//display("my name is ankita");/*this is multi line comment should be removed*/ 
input b; //inline comments//display("my name is ankita");/*this is multi line comment should be removed*/
endmodule

